LIBRARY ieee ;

USE ieee.std_logic_1164.all ;

PACKAGE fulladder_package IS
	COMPONENT fulladder
		PORT ( 
			Cin, A, B : IN STD_LOGIC ;
			S, Cout : OUT STD_LOGIC ) ;
	END COMPONENT ;
END fulladder_package ;
